module COMPUTE_BLOCK ( SET_TIME, ALARM, HRS, MINS, TOGGLE_SWITCH, CLK, RESETN,
                       DISPLAY, SPEAKER_OUT, TM_FIX );

input SET_TIME, ALARM, HRS, MINS, CLK, RESETN, TOGGLE_SWITCH, TM_FIX;
output SPEAKER_OUT;
output [10:0] DISPLAY;

wire TIM_AM_PM,ALM_AM_PM,KONNECT12;
wire [3:0] TIM_HRS,ALM_HRS;
wire [5:0] TIM_MINS,ALM_MINS;
reg INT_CLK;
wire [10:0] ALARM_BUS, TIME_BUS;

assign  DISPLAY = ALARM ? ALARM_BUS : TIME_BUS;

    CLOCK_GEN U7 ( .CLK(CLK), .RESETN(RESETN), .INT_CLK(INT_CLK) );

    TIME_BLOCK U1 ( .SET_TIME(SET_TIME), .HRS(HRS), .MINS(MINS),  
        .CLK(INT_CLK), .RESETN(RESETN), .ENABLE(!ALARM), 
        .HRS_OUT(TIM_HRS), .MINS_OUT(TIM_MINS), .AM_PM_OUT(TIM_AM_PM), 
        .DISPLAY_BUS(TIME_BUS) );

    ALARM_BLOCK  U2 ( .ALARM(ALARM), .HRS(HRS), .MINS(MINS), 
        .CLK(INT_CLK), .RESETN(RESETN), .ENABLE(ALARM),
        .HRS_OUT(ALM_HRS), .MINS_OUT(ALM_MINS), .AM_PM_OUT(ALM_AM_PM),
        .DISPLAY_BUS(ALARM_BUS) );

    COMPARATOR U4 ( .ALARM_HRS(ALM_HRS),.TIME_HRS(TIM_HRS), 
        .ALARM_MINS(ALM_MINS), .TIME_MINS(TIM_MINS),
        .ALARM_AM_PM(ALM_AM_PM), .TIME_AM_PM(TIM_AM_PM), .RINGER(KONNECT12) );

    ALARM_SM_2 U5 ( .COMPARE_IN(KONNECT12), .TOGGLE_ON(TOGGLE_SWITCH), 
        .CLOCK(INT_CLK), .RESETN(RESETN), .RING(SPEAKER_OUT) );

endmodule
